module BitSet(input [3:0]x,
			  input [1:0]index,
			  input value,
			  output [3:0]y);
	
endmodule